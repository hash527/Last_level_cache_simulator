package SnoopWrite;
    function automatic void SnoopedWrite(input_index,input_tag);
    // PASS
   endfunction
endpackage